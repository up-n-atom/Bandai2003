module BANDAI2003 (
    input CLK,
    input CEn,
    input WEn,
    input OEn,
    input SSn,
    output SO, /* Synchronous out */
    input RSTn,
    input [7:0] ADDR, /* A-1 to A3 + A15 to A18 */
    inout [7:0] DQ, /* Warning: Tri-state */
    output ROMCEn,
    output RAMCEn,
    output [9:0] RADDR /* ROM/RAM A15 to A24 - Starting at A-1 */
);

    reg [7:0] lckS; // Lock State - Addressed unlock sequence

    localparam ADDR_ACK = 8'h5A;
    localparam ADDR_NAK = 8'hA5;
    localparam ADDR_NIH = 8'hFF;

    wire LCKn = lckS != ADDR_NIH; // The end is nigh

    reg [17:0] shR; // Shift Register - Right

    // ¯\______/¯\_/¯\___/¯\_/¯\___/¯
    // Bit-stream - Invokes SYSTEM_CTRL1 (A0h) bit 7 to 1.
    localparam [17:0] bitS = {1'b0, 16'h28A0, 1'b0};

    assign SO = ~RSTn ? 1'bZ : shR[0]; // Change hi-Z on cart

    always @ (posedge CLK or negedge RSTn) begin
        if (~RSTn) begin
            shR <= {(18){1'b1}};
            lckS <= ADDR_ACK;
        end else if (LCKn && ADDR == lckS)
            case (ADDR)
                ADDR_ACK: lckS <= ADDR_NAK;
                ADDR_NAK: begin
                    shR <= bitS;
                    lckS <= ADDR_NIH;
                end
            endcase
        else
            shR <= {1'b1, shR[17:1]};
    end

    reg [7:0] laoR; // Linear Address Offset Register
    reg [9:0] bnkR [2:0]; // Bank Registers

    localparam ADDR_LAO = 8'hC0; // Linear Address Offset
    localparam ADDR_RAMB = 8'hC1; // RAM Bank
    localparam ADDR_ROMB0 = 8'hC2; // ROM Bank #0
    localparam ADDR_ROMB1 = 8'hC3; // ROM Bank #1
    localparam ADDR_RAMB_L = 8'hD0; // RAM Bank Low
    localparam ADDR_RAMB_H = 8'hD1; // RAM Bank High
    localparam ADDR_ROMB0_L = 8'hD2; // ROM Bank #0 Low
    localparam ADDR_ROMB0_H = 8'hD3; // ROM Bank #0 High
    localparam ADDR_ROMB1_L = 8'hD4; // ROM Bank #1 Low
    localparam ADDR_ROMB1_H = 8'hD5; // ROM Bank #1 High

    function [7:0] fDQ(
        input[7:0] ADDR
    );
        case (ADDR)
            ADDR_LAO: fDQ = laoR;
            ADDR_RAMB, ADDR_RAMB_L: fDQ = bnkR[0];
            ADDR_ROMB0, ADDR_ROMB0_L: fDQ = bnkR[1]
            ADDR_ROMB1, ADDR_ROMB1_L: fDQ = bnkR[2];
            ADDR_RAMB_H: fDQ = {6'b0, bnkR[0][9:8]};
            ADDR_ROMB0_H: fDQ = {6'b0, bnkR[1][9:8]};
            ADDR_ROMB1_H: fDQ = {6'b0, bnkR[2][9:8]};
            default: fDQ = 8'hFF;
        endcase
    endfunction

    wire seL = ~LCKn && ~(SSn & CEn);

    assign DQ = seL && ~OEn && WEn ? fDQ(ADDR) : 8'hZZ;
    wire [7:0] iDQ = DQ;

    wire rwC = OEn && WEn;

    integer i;

    always @(posedge rwC or negedge RSTn) begin
        if (~RSTn) begin
            laoR = 8'bFF;
            for (i = 0; i < 3; i = i + 1)
                bnkR[i] <= 10'h3FF;
        end else if (seL)
            case (ADDR)
                ADDR_LAO: laoR <= iDQ;
                ADDR_RAMB, ADDR_RAMB_L: bnkR[0] <= iDQ;
                ADDR_ROMB0, ADDR_ROMB0_L: bnkR[1] <= iDQ;
                ADDR_ROMB1, ADDR_ROMB1_L: bnkR[2] <= iDQ;
                ADDR_RAMB_H: bnkR[0][9:8] <= iDQ[1:0];
                ADDR_ROMB0_H: bnkR[1][9:8] <= iDQ[1:0];
                ADDR_ROMB1_H: bnkR[2][9:8] <= iDQ[1:0];
            endcase
    end

    wire rCE = ~LCKn && SSn && ~CEn;

    assign RAMCEn = ~(rCE && ADDR[7:4] == 4'h1);
    assign ROMCEn = ~(rCE && ADDR[7:4] > 4'h1);

    assign RADDR = ~RAMCEn || ~ROMCEn ? ADDR[7:4] > 4'h3 ? {laoR[5:0], ADDR[7:4]} : bnkR[ADDR[5:4] - 1] : 10'b0;

endmodule
